`timescale 1ns/1ps
module p1_tb;
    reg a, b, c, d;
    wire q;

    p1 uut (
        .a(a),
        .b(b),
        .c(c),
        .d(d),
        .q(q)
    );

    initial begin
        $monitor("a=%b , b=%b , c=%b , d=%b, q=%b", a, b, c, d, q);
        $dumpfile ("p1.vcd");
        $dumpvars (0,p1_tb);

        a = 0; b = 0; c = 0; d = 0; #10;
        a = 0; b = 0; c = 0; d = 1; #10;
        a = 0; b = 0; c = 1; d = 0; #10;
        a = 0; b = 0; c = 1; d = 1; #10;
        a = 0; b = 1; c = 0; d = 0; #10;
        a = 0; b = 1; c = 0; d = 1; #10;
        a = 1; b = 0; c = 0; d = 0; #10;
        a = 1; b = 0; c = 0; d = 1; #10;
        a = 1; b = 1; c = 0; d = 0; #10;
        a = 1; b = 1; c = 0; d = 1; #10;
        a = 1; b = 1; c = 1; d = 0; #10;
        a = 1; b = 1; c = 1; d = 1; #10;
        $finish;
    end
endmodule
