`timescale 1ps/1ps
module mux_8_1_tb;
    reg D1,D2,D3,D4,D5,D6,D7,D8,S1,S2,S3;
    wire q;  
    mux_8_1 uut(
    .D1(D1),
    .D2(D2),
    .D3(D3),
    .D4(D4),
    .D5(D5),
    .D6(D6),
    .D7(D7),
    .D8(D8),
    .S1(S1),
    .S2(S2),
    .S3(S3),
    .q(q)
    );
    initial begin 
        $dumpfile("mux_8_1.vcd");
        $dumpvars(0,mux_8_1_tb);

        S1=0; S2=0; S3=0; D1=1; D2=0; D3=0; D4=0; D5=0; D6=0; D7=0; D8=0; #10;
        S1=0; S2=0; S3=1; D1=0; D2=1; D3=0; D4=0; D5=0; D6=0; D7=0; D8=0; #10;
        S1=0; S2=1; S3=0; D1=0; D2=0; D3=1; D4=0; D5=0; D6=0; D7=0; D8=0; #10;
        S1=0; S2=1; S3=1; D1=0; D2=0; D3=0; D4=1; D5=0; D6=0; D7=0; D8=0; #10; 
        S1=1; S2=0; S3=0; D1=0; D2=0; D3=0; D4=0; D5=1; D6=0; D7=0; D8=0; #10;
        S1=1; S2=1; S3=1; D1=0; D2=0; D3=0; D4=0; D5=0; D6=1; D7=0; D8=0; #10;
        S1=1; S2=0; S3=0; D1=0; D2=0; D3=0; D4=0; D5=0; D6=0; D7=1; D8=0; #10;
        S1=1; S2=0; S3=1; D1=0; D2=0; D3=0; D4=0; D5=0; D6=0; D7=0; D8=1; #10;
        $finish;
    end
endmodule
